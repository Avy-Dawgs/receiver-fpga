/*
* Signal chain to measure power.
*/
module SignalChain
(
  input clk, 
  input rst, 
  input [11:0] data_i, 
  input valid_i,
  output data_o
); 

endmodule
