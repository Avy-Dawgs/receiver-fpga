/*
* Generates a sine wave at a particular frequency and sample rate.
*/
module SineGenerator
#(
  CLK_FREQ,
  FREQ,
  SAMP_RATE,
  DW
)
(
  input clk, 
  input rst, 
  input addr_i
); 

  
  

endmodule
